module logic_gates(
   input wire a,
   input wire b,
   output wire x
   );

assign x=a&b;
endmodule